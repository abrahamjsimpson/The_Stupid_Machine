
module OneBitProcessor
	(input clk,
	input reset,
	input en,
	input [1:0] inReg,
	output [6:0] outReg);


endmodule
	 